library ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

--library UNISIM;
--use UNISIM.VComponents.all;

package Config_LR is

end package Config_LR;



package body Config_LR is

end package body Config_LR;
